module top_module(output zero);
    
    assign zero = 0;

endmodule

//assign zero = 1'b0;
